module serial_buffer (
    input clock,
    input reset,
    
    input [31:0] addr_in,
    output reg [31:0] data_out,
    input re_in,
    input [31:0] data_in,
    input we_in,
    
    input s_data_valid_in, // Data to be read is available
    input [7:0] s_data_in, // Serial input data
    input s_data_ready_in, // Serial is ready to receive data
    output reg s_rden_out, // Serial read enable
    output reg [7:0] s_data_out, // Serial output data
    output reg s_wren_out // Serial write enable
);

    parameter MEM_ADDR = 16'hFFFF; // Memory-mapped address for the serial buffer

    // Read values (async)
    always @(*) begin
        case (addr_in[3:2])
            2'h0: data_out = {31'b0, s_data_valid_in}; // Status register: Data valid
            2'h1: data_out = {24'b0, s_data_in};       // Data register: Read data byte
            2'h2: data_out = {31'b0, s_data_ready_in}; // Ready register: Ready to receive
            2'h3: data_out = 32'b0;                   // Reserved or unused
            default: data_out = 32'b0;                // Default case for safety
        endcase
    end

    reg [7:0] sbyte; // Internal buffer for serial output data

    // Sequential logic for write and read enables
    always @(posedge clock or posedge reset) begin
        if (reset) begin
            s_rden_out <= 1'b0;
            s_wren_out <= 1'b0;
            sbyte <= 8'b0;
            s_data_out <= 8'b0; // Reset serial output
        end else begin
            s_rden_out <= 1'b0; // Default to no read operation
            s_wren_out <= 1'b0; // Default to no write operation

            // Check address and perform read/write operations
            if (addr_in[31:16] == MEM_ADDR) begin
                // Read operation: Triggered on read enable and correct address
                if (re_in && (addr_in[3:2] == 2'h1)) begin
                    s_rden_out <= 1'b1;
                end

                // Write operation: Triggered on write enable and correct address
                if (we_in && (addr_in[3:2] == 2'h3)) begin
                    sbyte <= data_in[7:0]; // Capture the lower byte of input data
                    s_data_out <= data_in[7:0]; // Procedural assignment to output
                    s_wren_out <= 1'b1;    // Assert write enable
                end
            end
        end
    end

endmodule
